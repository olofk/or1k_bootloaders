@00000000
18000000
18609100
18800000
9C8000FF
D8032000
D8032001
18E0000F
A8E74240
18800000
9C800080
D8032000
B8840041
18C00000
9CC60001
E4063800
0FFFFFFE
15000000
E4040000
15000000
0FFFFFF7
15000000
03FFFFF3
15000000
